`timescale 1ns/1ns

module Q6_myBarrelVectorCondition (output [15:0]W, input [15:0]D, [15:0]N);
	wire [15:0]XV = 0;

	assign #(317) W = N[0]?{D[15:0]}:
			N[1]?{XV[0:0], D[15:1]}:
			N[2]?{XV[1:0], D[15:2]}:
			N[3]?{XV[2:0], D[15:3]}:
			N[4]?{XV[3:0], D[15:4]}:
			N[5]?{XV[4:0], D[15:5]}:
			N[6]?{XV[5:0], D[15:6]}:
			N[7]?{XV[6:0], D[15:7]}:
			N[8]?{XV[7:0], D[15:8]}:
			N[9]?{XV[8:0], D[15:9]}:
			N[10]?{XV[9:0], D[15:10]}:
			N[11]?{XV[10:0], D[15:11]}:
			N[12]?{XV[11:0], D[15:12]}:
			N[13]?{XV[12:0], D[15:13]}:
			N[14]?{XV[13:0], D[15:14]}:
			N[15]?{XV[14:0], D[15:15]}:XV[15:0];
endmodule