`timescale 1ns/1ns

module Q8_myBarrelNmos(output [7:0]W, input [7:0]D,  [7:0]N);	
	supply0 Gnd;
	nmos#(3,4,5) (W[0], D[0], N[0]), (W[0], D[1], N[1]), (W[0], D[2], N[2]), (W[0], D[3], N[3]), (W[0], D[4], N[4]), (W[0], D[5], N[5]), (W[0], D[6], N[6]), (W[0], D[7], N[7]); 
	nmos#(3,4,5) (W[1], D[1], N[0]), (W[1], D[2], N[1]), (W[1], D[3], N[2]), (W[1], D[4], N[3]), (W[1], D[5], N[4]), (W[1], D[6], N[5]), (W[1], D[7], N[6]), (W[1], Gnd, N[7]); 
	nmos#(3,4,5) (W[2], D[2], N[0]), (W[2], D[3], N[1]), (W[2], D[4], N[2]), (W[2], D[5], N[3]), (W[2], D[6], N[4]), (W[2], D[7], N[5]), (W[2], Gnd, N[6]), (W[2], Gnd, N[7]); 
	nmos#(3,4,5) (W[3], D[3], N[0]), (W[3], D[4], N[1]), (W[3], D[5], N[2]), (W[3], D[6], N[3]), (W[3], D[7], N[4]), (W[3], Gnd, N[5]), (W[3], Gnd, N[6]), (W[3], Gnd, N[7]); 
	nmos#(3,4,5) (W[4], D[4], N[0]), (W[4], D[5], N[1]), (W[4], D[6], N[2]), (W[4], D[7], N[3]), (W[4], Gnd, N[4]), (W[4], Gnd, N[5]), (W[4], Gnd, N[6]), (W[4], Gnd, N[7]); 
	nmos#(3,4,5) (W[5], D[5], N[0]), (W[5], D[6], N[1]), (W[5], D[7], N[2]), (W[5], Gnd, N[3]), (W[5], Gnd, N[4]), (W[5], Gnd, N[5]), (W[5], Gnd, N[6]), (W[5], Gnd, N[7]); 
	nmos#(3,4,5) (W[6], D[6], N[0]), (W[6], D[7], N[1]), (W[6], Gnd, N[2]), (W[6], Gnd, N[3]), (W[6], Gnd, N[4]), (W[6], Gnd, N[5]), (W[6], Gnd, N[6]), (W[6], Gnd, N[7]); 
	nmos#(3,4,5) (W[7], D[7], N[0]), (W[7], Gnd, N[1]), (W[7], Gnd, N[2]), (W[7], Gnd, N[3]), (W[7], Gnd, N[4]), (W[7], Gnd, N[5]), (W[7], Gnd, N[6]), (W[7], Gnd, N[7]);
endmodule